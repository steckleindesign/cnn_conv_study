`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 01/10/2025 03:15:37 PM
// Design Name: 
// Module Name: windowed_feature
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module windowed_feature #(parameter LAST_COL = 0) (
    input  in0,
    input  in1,
    output feature
);

    

endmodule
